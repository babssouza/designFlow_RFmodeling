.SUBCKT		tstFixture_S2-LP_081920_085345_10016
+			Port1_1
+			Port1_3
+			Port2_5
+			Port2_7
*The following is the Cadence MCP(model connection protocol) Section
***********************************
*[MCP Begin]
*[MCP Ver] 1.1
*[MCP Source] Cadence Design Systems, Inc. PowerSI 16.0.0.02091.0   000 8/19/2020
*
***********************************
*
*[REM]The following is the info for non-circuit ports
*[REM]**********************************
*[Connection] general unnamed 8
*[Power Nets]
*[Ground Nets]
*Port1_N_3	Port1_3	GND	0.1758930	0.0640180
*Port1_N_4	Port1_3	GND	0.1758930	0.1140180
*Port2_N_7	Port2_7	GND	0.2701780	0.1140180
*Port2_N_8	Port2_7	GND	0.2231330	0.0640580
*[Signal Nets]
*Port1_P_1	Port1_1	TX	0.1772270	0.0640010
*Port1_P_2	Port1_1	TX	0.1772270	0.1140010
*Port2_P_5	Port2_5	TX	0.2221300	0.0639980
*Port2_P_6	Port2_5	TX	0.2686770	0.1140010
*
*[MCP End]
*
*This concludes the MCP section
*Define the S element, the Model file is output from BNP

.MODEL   Spara   S		
+		BNPFILE = "tstFixture_S2-LP_081920_085345_10016.bnp"

S		
+			Port1_1	Port1_3
+			Port2_5	Port2_7
+			MNAME = Spara

*
.ENDS
*
*
