.SUBCKT		tstFixture_S2-LP_081920_102238_10016
+			Port1_1
+			Port1_3
*The following is the Cadence MCP(model connection protocol) Section
***********************************
*[MCP Begin]
*[MCP Ver] 1.1
*[MCP Source] Cadence Design Systems, Inc. PowerSI 16.0.0.02091.0   000 8/19/2020
*
***********************************
*
*[REM]The following is the info for non-circuit ports
*[REM]**********************************
*[Connection] general unnamed 4
*[Power Nets]
*[Ground Nets]
*Port1_N_3	Port1_3	GND	0.2703590	0.1605600
*Port1_N_4	Port1_3	GND	0.1760740	0.1605600
*[Signal Nets]
*Port1_P_1	Port1_1	TX	0.2688580	0.1605430
*Port1_P_2	Port1_1	TX	0.1774080	0.1605430
*
*[MCP End]
*
*This concludes the MCP section
*Define the S element, the Model file is output from BNP

.MODEL   Spara   S		
+		BNPFILE = "tstFixture_S2-LP_081920_102238_10016.bnp"

S		
+			Port1_1	Port1_3
+			MNAME = Spara

*
.ENDS
*
*
